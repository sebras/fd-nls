HELP.TXT

Hj�lp:

Detta program spelar in filpositionsinformation f�r eventuellt �terskapande
via UNFORMAT.

Syntax:

MIRROR [enhet:]
MIRROR [/PARTN]

  /PARTN    Lagrar en s�kerhetskopia av partitionstabellerna i en PARNSAV.FIL
              p� disketten i A:-enheten. Partitionstabellerna kan �terskapas
	      med UNFORMAT version 0.8.





